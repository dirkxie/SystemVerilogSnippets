module FIFO_async
