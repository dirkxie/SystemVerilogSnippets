module GrayCounter
# (
 parameter COUNTER_WIDTH = 4)
